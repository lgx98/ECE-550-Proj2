module regfile (clock,
                ctrl_writeEnable,
                ctrl_reset,
                ctrl_writeReg,
                ctrl_readRegA,
                ctrl_readRegB,
                data_writeReg,
                data_readRegA,
                data_readRegB);
    
    input clock, ctrl_writeEnable, ctrl_reset;
    input [4:0] ctrl_writeReg, ctrl_readRegA, ctrl_readRegB;
    input [31:0] data_writeReg;
    
    output [31:0] data_readRegA, data_readRegB;
    
    /* YOUR CODE HERE */
    
endmodule
